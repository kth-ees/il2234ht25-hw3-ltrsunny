module sequence_detector_structural (
    input logic clk,
    input logic rst_n,
    input logic input_sequence,
    output logic detected
);

	// …
	// Add your description here
	// …

endmodule

