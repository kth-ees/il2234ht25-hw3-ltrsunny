module sequence_detector_behavioral (
    input logic clk,
    input logic rst_n,
    input logic input_sequence,
    output logic detected
);

	// …
	// Add your description here
	// …

endmodule