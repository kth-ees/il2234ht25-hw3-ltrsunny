module serial_communication(
    input logic clk,
    input logic rst_n,
    input logic serData,
    output logic outValid
);

	// …
	// Add your description here
	// …


endmodule