module conversion_system_mealy (
    input logic clk,
    input logic rst_n,
    input logic x,
    output logic z
);

	// …
	// Add your description here
	// …


endmodule