module sin (
    input  logic        clk,
    input  logic        rst_n,
    input  logic [15:0] x,
    input  logic        start,
    output logic [15:0] result,
    output logic        done
);

	// …
	// Add your description here
	// …

endmodule