module conversion_system_moore (
    input logic clk,
    input logic rst_n,
    input logic x,
    output logic z
);

	// …
	// Add your description here
	// …

endmodule
