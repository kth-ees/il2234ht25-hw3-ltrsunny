module average_calc_controller #(parameter n = 4) (
    input logic clk,
    input logic rst_n,
    input logic start,
    output logic init_sum,
    output logic init_shift,
    output logic load,
    output logic shift,
    output logic done
);

	// …
	// Add your description here
	// …

endmodule